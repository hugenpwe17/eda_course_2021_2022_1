module h_adder1(
	input ain,
	input bin,
	
	output sout,
	output cout
	);
	// reg
	
	// wire
	
	// main code
	assign sout = ain ^ bin;
	assign cout = ain & bin;

endmodule