library verilog;
use verilog.vl_types.all;
entity main_vlg_check_tst is
    port(
        clk_div         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end main_vlg_check_tst;
