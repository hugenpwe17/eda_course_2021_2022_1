// key_led
module key_led(
	input sys_clk,
	input sys_rst_n,
	input [3:0] key,
	
	output reg [3:0] led);
	
	//reg
	reg [23:0] cnt;
	reg [1:0] led_ctl;
	
	// 0.2s conter
	always@(posedge sys_clk, negedge sys_rst_n)begin
		if(!sys_rst_n) 
			cnt <= 24'd9_999_999;
		else if(cnt <= 24'd9_999_999)
			cnt <= cnt + 1;
		else
			cnt <= 0;
	end
	
	// led status select
	always@(posedge sys_clk, negedge sys_rst_n)begin
		if(!sys_rst_n)
			led_ctl <= 2'b00;
		else if(cnt == 24'd9_999_999)
			led_ctl <= led_ctl + 1'b1;
		else
			led_ctl <= led_ctl;
	end
	
	// detect key
	always@(posedge sys_clk, negedge sys_rst_n)begin
		if(!sys_rst_n)
			led <= 4'b0000;
		else if(key[0] == 0)
			case(led_ctl)
				2'b00 : led <= 4'b1000;
				2'b01 : led <= 4'b0100;
				2'b10 : led <= 4'b0010;
				2'b11 : led <= 4'b0001;
				default : led <= 4'b0000;
			endcase
		else if(key[1] == 0)
			case(led_ctl)
				2'b00 : led <= 4'b0001;
				2'b01 : led <= 4'b0010;
				2'b10 : led <= 4'b0100;
				2'b11 : led <= 4'b1000;
				default : led <= 4'b0000;
			endcase
		else if(key[2] == 0)
			case(led_ctl)
				2'b00 : led <= 4'b1010;
				2'b01 : led <= 4'b0101;
				2'b10 : led <= 4'b1010;
				2'b11 : led <= 4'b0101;
				default : led <= 4'b0000;
			endcase
		else if(key[3] == 0)
			led = 4'b1111;
		else
			led <= 4'b0000;
			//case(led_ctl)
			//	2'b00 : led <= 4'b1000;
			//	2'b01 : led <= 4'b0000;
			//	2'b10 : led <= 4'b1000;
			//	2'b11 : led <= 4'b0000;
			//	default : led <= 4'b0000;
			//endcase
	end
	
endmodule