module cnt_hex_seg_dync_top (
    input clk,
    input rst_n,

    output [7:0] seg,
    output [2:0] sel
);
    
endmodule